.title KiCad schematic
.include "models/C2012C0G2A102J060AA_p.mod"
.include "models/C2012X7R2A104K125AA_p.mod"
.include "models/CGJ4C2C0G2A101J060AA_p.mod"
.include "models/MBRS340T3.LIB"
.include "models/PCF1C101MCL1GS_v100.lib"
.include "models/PCV1J220MCL6GS_v100.lib"
.include "models/SML-D12P8W.lib"
.include "models/ZXMP7A17K.lib"
.include "models/lm3485.lib"
XU5 /SENSE 0 /FB /ADJ /PGATE VCC LM3485
R1 VCC /ADJ 24.0k
XU2 VCC /ADJ C2012C0G2A102J060AA_p
XU3 VCC 0 C2012X7R2A104K125AA_p
XU7 /SENSE /PGATE VCC ZXMP7A17K
XU6 /OUT /FB CGJ4C2C0G2A101J060AA_p
L1 /SENSE /OUT 22u rser=0.028
R2 /OUT /FB {Rfb}
R3 /FB 0 {Rref}
XU8 /COUT 0 PCF1C101MCL1GS
XU1 VCC 0 PCV1J220MCL6GS
R5 /OUT /PWRON 562
D2 /PWRON 0 SML-D12P8W
R4 /OUT /COUT {Rser_Cout}
XU4 VCC 0 C2012X7R2A104K125AA_p
D1 0 /SENSE Dmbrs340
V1 VCC 0 {VIN}
I1 /OUT 0 {ILOAD}
.end
